library verilog;
use verilog.vl_types.all;
entity ex1_tb is
end ex1_tb;
