library verilog;
use verilog.vl_types.all;
entity c1_tb is
end c1_tb;
