library verilog;
use verilog.vl_types.all;
entity counter_tb is
    generic(
        size            : integer := 8
    );
end counter_tb;
