library verilog;
use verilog.vl_types.all;
entity ex1b_tb is
end ex1b_tb;
