library verilog;
use verilog.vl_types.all;
entity dff_tb is
end dff_tb;
