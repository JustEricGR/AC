library verilog;
use verilog.vl_types.all;
entity ex1b is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        f2              : out    vl_logic
    );
end ex1b;
