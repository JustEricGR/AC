module main ;
  initial
  $display(" H e l l o , w o r l d ! ") ;
endmodule