library verilog;
use verilog.vl_types.all;
entity sha2indpath_tb is
end sha2indpath_tb;
