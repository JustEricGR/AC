library verilog;
use verilog.vl_types.all;
entity regfl_tb is
end regfl_tb;
